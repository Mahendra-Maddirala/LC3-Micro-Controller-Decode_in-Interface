//decode_test_pkg
package decode_test_pkg;
  import uvm_pkg::*;
  import decode_in_pkg::*;

  `include "uvm_macros.svh"
  `include "test_top.sv"

endpackage: decode_test_pkg
